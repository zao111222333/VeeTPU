`timescale 1ns/1ps
module top_tb();
parameter clk_period = 2;
reg clk;
reg [1:0] mode_sel;
reg rstn;

initial begin
    rstn <= 0;
	 clk  <= 0;
	 #clk_period rstn <= 1'b1;
end

initial begin
 forever #(clk_period/2) clk <= ~clk; 
end

reg [15:0] a[15:0];
reg [15:0] b[15:0];

initial begin
    $dumpfile("wave.vcd");
    $dumpvars(0,top_tb);
end
//FP32 test
initial begin
    a[ 0]<=16'b0;
    a[ 1]<=16'b0;
    a[ 2]<=16'b0;
    a[ 3]<=16'b0;
    a[ 4]<=16'b0;
    a[ 5]<=16'b0;
    a[ 6]<=16'b0;
    a[ 7]<=16'b0;
    a[ 8]<=16'b0;
    a[ 9]<=16'b0;
    a[10]<=16'b0;
    a[11]<=16'b0;
    a[12]<=16'b0;
    a[13]<=16'b0;
    a[14]<=16'b0;
    a[15]<=16'b0;
    b[ 0]<=16'b0;
    b[ 1]<=16'b0;
    b[ 2]<=16'b0;
    b[ 3]<=16'b0;
    b[ 4]<=16'b0;
    b[ 5]<=16'b0;
    b[ 6]<=16'b0;
    b[ 7]<=16'b0;
    b[ 8]<=16'b0;
    b[ 9]<=16'b0;
    b[10]<=16'b0;
    b[11]<=16'b0;
    b[12]<=16'b0;
    b[13]<=16'b0;
    b[14]<=16'b0;
    b[15]<=16'b0;
#(clk_period+clk_period/2)
    a[ 0]<=16'b0_10001_1010000000;
    a[ 1]<=16'b0_10100_0101001000;
    a[ 2]<=16'b0_10111_1010011010;
    a[ 3]<=16'b0_10001_0111100000;
    a[ 4]<=16'b0_10001_0100000100;
    a[ 5]<=16'b0_10001_0100000010;
    a[ 6]<=16'b0_10001_0100000001;
    a[ 7]<=16'b0_10001_1000000010;
    a[ 8]<=16'b0_10001_1010000000;
    a[ 9]<=16'b0_10000_1000000000;
    a[10]<=16'b0_10000_0100000100;
    a[11]<=16'b0_10000_0100000010;
    a[12]<=16'b0_10000_0100000001;
    a[13]<=16'b0_10000_1000000010;
    a[14]<=16'b0_10000_1010000000;
    a[15]<=16'b0_10000_1000000000;
    b[ 0]<=16'b0_10000_0100000000;
    b[ 1]<=16'b0_10000_0111100000;
    b[ 2]<=16'b0_10000_0100000100;
    b[ 3]<=16'b0_10000_0100000010;
    b[ 4]<=16'b0_10000_0100000001;
    b[ 5]<=16'b0_10000_1000000010;
    b[ 6]<=16'b0_10000_0100000100;
    b[ 7]<=16'b0_10000_0100000010;
    b[ 8]<=16'b0_10000_0100000001;
    b[ 9]<=16'b0_10000_1000000010;
    b[10]<=16'b0_10000_0100000001;
    b[11]<=16'b0_10000_1000000010;
    b[12]<=16'b0_10000_0100000100;
    b[13]<=16'b0_10000_0100000010;
    b[14]<=16'b0_10000_0100000001;
    b[15]<=16'b0_10000_1000000010;
#clk_period
    a[ 0]<=16'b0_10000_1000000000;
    a[ 1]<=16'b0_10000_1000000000;
    a[ 2]<=16'b0_10000_1000000000;
    a[ 3]<=16'b0_10000_1000000000;
    a[ 4]<=16'b0_10000_1000000000;
    a[ 5]<=16'b0_10000_1000000000;
    a[ 6]<=16'b0_10000_1000000000;
    a[ 7]<=16'b0_10000_1000000000;
    a[ 8]<=16'b0_10000_1000000000;
    a[ 9]<=16'b0_10000_1000000000;
    a[10]<=16'b0_10000_1000000000;
    a[11]<=16'b0_10000_1000000000;
    a[12]<=16'b0_10000_1000000000;
    a[13]<=16'b0_10000_1000000000;
    a[14]<=16'b0_10000_1000000000;
    a[15]<=16'b0_10000_1000000000;
    b[ 0]<=16'b0_01111_0000000000;
    b[ 1]<=16'b0_01111_0000000000;
    b[ 2]<=16'b0_01111_0000000000;
    b[ 3]<=16'b0_01111_0000000000;
    b[ 4]<=16'b0_01111_0000000000;
    b[ 5]<=16'b0_01111_0000000000;
    b[ 6]<=16'b0_01111_0000000000;
    b[ 7]<=16'b0_01111_0000000000;
    b[ 8]<=16'b0_10000_1000000000;
    b[ 9]<=16'b0_10000_1000000000;
    b[10]<=16'b0_10000_1000000000;
    b[11]<=16'b0_10000_1000000000;
    b[12]<=16'b0_10000_1000000000;
    b[13]<=16'b0_10000_1000000000;
    b[14]<=16'b0_10000_1000000000;
    b[15]<=16'b0_10000_1000000000;
#clk_period
    a[ 0]<=16'b0;
    a[ 1]<=16'b0;
    a[ 2]<=16'b0;
    a[ 3]<=16'b0;
    a[ 4]<=16'b0;
    a[ 5]<=16'b0;
    a[ 6]<=16'b0;
    a[ 7]<=16'b0;
    a[ 8]<=16'b0;
    a[ 9]<=16'b0;
    a[10]<=16'b0;
    a[11]<=16'b0;
    a[12]<=16'b0;
    a[13]<=16'b0;
    a[14]<=16'b0;
    a[15]<=16'b0;
    b[ 0]<=16'b0;
    b[ 1]<=16'b0;
    b[ 2]<=16'b0;
    b[ 3]<=16'b0;
    b[ 4]<=16'b0;
    b[ 5]<=16'b0;
    b[ 6]<=16'b0;
    b[ 7]<=16'b0;
    b[ 8]<=16'b0;
    b[ 9]<=16'b0;
    b[10]<=16'b0;
    b[11]<=16'b0;
    b[12]<=16'b0;
    b[13]<=16'b0;
    b[14]<=16'b0;
    b[15]<=16'b0;
end

/*FP16 test
initial begin
    a[ 0]<=16'b0;
    a[ 1]<=16'b0;
    a[ 2]<=16'b0;
    a[ 3]<=16'b0;
    a[ 4]<=16'b0;
    a[ 5]<=16'b0;
    a[ 6]<=16'b0;
    a[ 7]<=16'b0;
    a[ 8]<=16'b0;
    a[ 9]<=16'b0;
    a[10]<=16'b0;
    a[11]<=16'b0;
    a[12]<=16'b0;
    a[13]<=16'b0;
    a[14]<=16'b0;
    a[15]<=16'b0;
    b[ 0]<=16'b0;
    b[ 1]<=16'b0;
    b[ 2]<=16'b0;
    b[ 3]<=16'b0;
    b[ 4]<=16'b0;
    b[ 5]<=16'b0;
    b[ 6]<=16'b0;
    b[ 7]<=16'b0;
    b[ 8]<=16'b0;
    b[ 9]<=16'b0;
    b[10]<=16'b0;
    b[11]<=16'b0;
    b[12]<=16'b0;
    b[13]<=16'b0;
    b[14]<=16'b0;
    b[15]<=16'b0;
#(clk_period+clk_period/2)
    a[ 0] <= 16'b0_10001_1010000000;
    a[ 1] <= 16'b0_10100_0101001000;
    a[ 2] <= 16'b0_10011_1010011010;
    a[ 3] <= 16'b0_10001_0111100000;
    a[ 4] <= 16'b0_10001_0100000100;
    a[ 5] <= 16'b0_10001_0100000010;
    a[ 6] <= 16'b0_10001_0100000001;
    a[ 7] <= 16'b0_10001_1000000010;
    a[ 8] <= 16'b0_10001_1010000000;
    a[ 9] <= 16'b0_10001_1000000000;
    a[10] <= 16'b0_10001_0100000100;
    a[11] <= 16'b0_10001_0100000010;
    a[12] <= 16'b0_10001_0100000001;
    a[13] <= 16'b0_10001_1000000010;
    a[14] <= 16'b0_10001_1010000000;
    a[15] <= 16'b0_10001_1000000000;
    
    b[ 0] <= 16'b0_10001_0100000000;
    b[ 1] <= 16'b0_10001_0111100000;
    b[ 2] <= 16'b0_10001_0100000100;
    b[ 3] <= 16'b0_10001_0100000010;
    b[ 4] <= 16'b0_10001_0100000001;
    b[ 5] <= 16'b0_10001_1000000010;
    b[ 6] <= 16'b0_10001_0100000100;
    b[ 7] <= 16'b0_10001_0100000010;
    b[ 8] <= 16'b0_10001_0100000001;
    b[ 9] <= 16'b0_10001_1000000010;
    b[10] <= 16'b0_10001_0100000001;
    b[11] <= 16'b0_10001_1000000010;
    b[12] <= 16'b0_10001_0100000100;
    b[13] <= 16'b0_10001_0100000010;
    b[14] <= 16'b0_10001_0100000001;
    b[15] <= 16'b0_10001_1000000010;
#clk_period
    a[ 0]<=16'b0_10000_1000000000;
    a[ 1]<=16'b0_10000_1000000000;
    a[ 2]<=16'b0_10000_1000000000;
    a[ 3]<=16'b0_10000_1000000000;
    a[ 4]<=16'b0_10000_1000000000;
    a[ 5]<=16'b0_10000_1000000000;
    a[ 6]<=16'b0_10000_1000000000;
    a[ 7]<=16'b0_10000_1000000000;
    a[ 8]<=16'b0_10000_1000000000;
    a[ 9]<=16'b0_10000_1000000000;
    a[10]<=16'b0_10000_1000000000;
    a[11]<=16'b0_10000_1000000000;
    a[12]<=16'b0_10000_1000000000;
    a[13]<=16'b0_10000_1000000000;
    a[14]<=16'b0_10000_1000000000;
    a[15]<=16'b0_10000_1000000000;
    b[ 0]<=16'b0_10000_1000000000;
    b[ 1]<=16'b0_10000_1000000000;
    b[ 2]<=16'b0_10000_1000000000;
    b[ 3]<=16'b0_10000_1000000000;
    b[ 4]<=16'b0_10000_1000000000;
    b[ 5]<=16'b0_10000_1000000000;
    b[ 6]<=16'b0_10000_1000000000;
    b[ 7]<=16'b0_10000_1000000000;
    b[ 8]<=16'b0_10000_1000000000;
    b[ 9]<=16'b0_10000_1000000000;
    b[10]<=16'b0_10000_1000000000;
    b[11]<=16'b0_10000_1000000000;
    b[12]<=16'b0_10000_1000000000;
    b[13]<=16'b0_10000_1000000000;
    b[14]<=16'b0_10000_1000000000;
    b[15]<=16'b0_10000_1000000000;
#clk_period
    a[ 0]<=16'b0;
    a[ 1]<=16'b0;
    a[ 2]<=16'b0;
    a[ 3]<=16'b0;
    a[ 4]<=16'b0;
    a[ 5]<=16'b0;
    a[ 6]<=16'b0;
    a[ 7]<=16'b0;
    a[ 8]<=16'b0;
    a[ 9]<=16'b0;
    a[10]<=16'b0;
    a[11]<=16'b0;
    a[12]<=16'b0;
    a[13]<=16'b0;
    a[14]<=16'b0;
    a[15]<=16'b0;
    b[ 0]<=16'b0;
    b[ 1]<=16'b0;
    b[ 2]<=16'b0;
    b[ 3]<=16'b0;
    b[ 4]<=16'b0;
    b[ 5]<=16'b0;
    b[ 6]<=16'b0;
    b[ 7]<=16'b0;
    b[ 8]<=16'b0;
    b[ 9]<=16'b0;
    b[10]<=16'b0;
    b[11]<=16'b0;
    b[12]<=16'b0;
    b[13]<=16'b0;
    b[14]<=16'b0;
    b[15]<=16'b0;
end
*/

wire [63:0] r;
wire out_en;
PE_16in_top u_test(
    .clk(clk),
    .rstn(rstn),
    .mode_sel(2'b01),
    .A({a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15]}),
    .B({b[0],b[1],b[2],b[3],b[4],b[5],b[6],b[7],b[8],b[9],b[10],b[11],b[12],b[13],b[14],b[15]}),
    .acc_num(3),
    .result(r),
    .out_en(out_en)
    );
/*
integer out_file;

initial
begin
    out_file = $fopen("./out_put_file.txt","w");
end
initial
begin
#12
    $fwrite(out_file,"%h",r);
#2
    $fwrite(out_file,"%h",r);
#2  $finish;
end
*/
endmodule
